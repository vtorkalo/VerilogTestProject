module lcd_module(
  input logic CLK,
  input logic RESET,
  input logic sendText,
  input logic [8 * LINE_LENGTH : 1] line1,
  input logic [8 * LINE_LENGTH : 1] line2,
  inout [3:0] LCD_D,
  output logic LCD_RS,
  output logic LCD_E,
  output logic LCD_RW,
  output logic sendingDone
);

localparam LINE_LENGTH = 6'd16;

always_ff @(posedge CLK, posedge RESET)
begin
   if (RESET)
   begin
      state_reg <= not_init;
   end
   else
   begin
      state_reg <= state_next;
   end
end

typedef enum bit[4:0] {not_init, send_init_command, init_done, send_text, sending_done, idle} state_type;
state_type state_reg, state_next;


always_comb
begin
   state_next = state_reg;
   startInit_tick = 1'b0;
   sendText_tick = 1'b0;

     
   case (state_reg)
      not_init:
      begin
        if (sendText)
           state_next = send_init_command;
      end
      send_init_command:
      begin
         startInit_tick = 1'b1;      
         if (initDone)
            state_next = init_done;
      end
      init_done:
      begin
         state_next = send_text;
      end      
      send_text:
      begin
         sendText_tick = 1'b1;
         if (sendingDone)
            state_next = idle;
      end
      idle:
      begin
        if (sendText)
        begin
           state_next = send_text;
        end 
      end
   endcase

end

logic startInit_tick;
logic initDone;

logic LCD_D_IN_init; 
logic [3:0] LCD_D_init;
logic LCD_E_init;
logic LCD_RW_init;
logic LCD_RS_init;
logic READ_init;

logic LCD_D_IN_text;
logic [3:0] LCD_D_text;
logic LCD_E_text;
logic LCD_RW_text;
logic LCD_RS_text;
logic READ_text;


logic notInitialized;
assign notInitialized = state_reg == not_init | state_reg == send_init_command;

assign LCD_D = notInitialized ? (READ_init ? 4'bZZZZ : LCD_D_init)
                              : (READ_text ? 4'bZZZZ : LCD_D_text);
                              
assign busy_flag_init =  LCD_D[3];
assign busy_flag_text = LCD_D[3];

assign LCD_E = notInitialized ? LCD_E_init : LCD_E_text;
assign LCD_RW = notInitialized ? LCD_RW_init : LCD_RW_text;
assign LCD_RS = notInitialized ? LCD_RS_init : LCD_RS_text;



lcd_init lcd_init(.CLK(CLK),
   .RESET(RESET),
   .startInit(startInit_tick),
   .LCD_D(LCD_D_init),
   .busy_flag(busy_flag_init),
   .LCD_E(LCD_E_init),
   .LCD_RW(LCD_RW_init),
   .LCD_RS(LCD_RS_init),
   .initDone(initDone),
   .READ(READ_init));

logic sendText_tick;


lcd_send_text lcd_text(.CLK(CLK),
   .RESET(RESET),
   .sendText(sendText_tick),
   .line1(line1),
   .line2(line2),
   .LCD_D(LCD_D_text),
   .busy_flag(busy_flag_text),
   .LCD_E(LCD_E_text),
   .LCD_RW(LCD_RW_text),
   .LCD_RS(LCD_RS_text),
   .READ(READ_text),
   .sendingDone(sendingDone));
   
   
endmodule